// =====================================
//Simulation model of SRAM
//Author:     HuRui
//Modules:    sim_ram
//assume legal address
//=====================================

module sim_ram#(
    parameter DP = 512,//depth
    parameter DW = 32,//data width
    parameter MW= 4,//mask width
    parameter AW = 32,//address width
    parameter FORCE_X2ZERO = 0,
    parameter ITCM = 0,//instantiate as ITCM RAM
    parameter DTCM = 0 //instantiate as DTCM RAM
) (
    input  clk,
    input[DW-1:0] din,
    input[AW-1:0] addr,
    input we,
    input[MW-1:0] wem,//write enable mask
    output[DW-1:0] dout
);

    reg [DW-1:0] mem_r[0:DP-1];
    reg [AW-1:0] addr_r;
    wire [MW-1:0] wen;
    wire ren;

    assign ren = ~we;
    assign wen = ({MW{we}} & wem);

    //the output will holdup
    always @(posedge clk ) begin
        if(ren) begin
            addr_r <= addr;
        end
    end
<<<<<<< HEAD
    
    wire[DW-1:0] dout_pre;
    assign dout_pre = mem_r[addr];
    assign dout = dout_pre;
    
   
    initial begin
        if (ITCM==1) begin
            mem_r[0] = 32'b0000000_00000_00000_001_00001_011_0111;//lui
            mem_r[1] = 32'b0000000_00000_00000_001_00001_011_0110;//lui
            mem_r[2] = 32'b0000000_00000_00000_001_00001_011_0101;//lui
            mem_r[3] = 32'b0000000_00000_00000_001_00001_011_0100;//lui
=======
    
    genvar i;
    generate
        for(i = 0; i<MW; i = i + 1) begin
            if((8*i+8) > DW) begin
                always @(posedge clk) begin
                    if (wen[i]) begin
                        mem_r[addr][DW-1:8*i] <= din[DW-1:8*i];
                    end
                end
            end
            else begin
                always @(posedge clk) begin
                    if (wen[i]) begin
                        mem_r[addr][8*i+7:8*i] <= din[8*i+7:8*i];
                    end
                end
            end
        end
    endgenerate
    
    wire [DW-1:0] dout_pre;
    assign dout_pre = mem_r[addr_r];
    assign dout = dout_pre;
    /*
      generate
       if(FORCE_X2ZERO == 1) begin: force_x_to_zero
          for (i = 0; i < DW; i = i+1) begin:force_x_gen 
              `ifndef SYNTHESIS//{
             assign dout[i] = (dout_pre[i] === 1'bx) ? 1'b0 : dout_pre[i];
              `else//}{
             assign dout[i] = dout_pre[i];
              `endif//}
          end
       end
       else begin:no_force_x_to_zero
         assign dout = dout_pre;
       end
      endgenerate
    */
    
    
    initial begin
        if (ITCM == 1) begin
            mem_r[0] <= 32'b0000000_00000_00000_001_00001_011_0111;//lui
            mem_r[1] <= 32'b0000000_00000_00000_001_00001_011_0111;//lui
            mem_r[2] <= 32'b0000000_00000_00000_001_00001_011_0111;//lui
            mem_r[3] <= 32'b0000000_00000_00000_001_00001_011_0111;//lui
>>>>>>> 3cc96cc598ee1870011e45f9ad3faf27b1a26f50
        end
    end

endmodule
