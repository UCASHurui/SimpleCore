module exu_regfile (
    
);
    
endmodule